`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/07 13:14:01
// Design Name: 
// Module Name: SPI_Master
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SPI_Master (
    // Global Signals
    input logic clk,
    input logic reset,
    // Internal Signals
    input logic start,
    input logic [7:0] tx_data,
    output logic [7:0] rx_data,
    output logic tx_ready,
    output logic done,
    // External SPI Signals
    output logic SCLK,
    output logic MOSI,
    input logic MISO
    // Slave Select�� �Ϲ������� GPIO ������ ����ǰ�, ���� wrapper ��⿡�� ����.
);


    // ���� ���迡����, SCLK�� ���ֱ⸦ CPO(SCLK=0), ������ �� �ֱ⸦ CP1(SCLK=1)�� �����ϰ�,
    // �� State���� MOSI, MISO ��ȣ�� ó���ϴ� ������� ����.
    typedef enum {
        IDLE,
        CP0,
        CP1
    } state_t;

    state_t c_state, n_state;

    logic [7:0] tx_data_reg, tx_data_next;          // To prevent Latch
    logic [7:0] rx_data_reg, rx_data_next;          // To prevent Latch

    logic [5:0] sclk_count_reg, sclk_count_next;    // To prevent Latch
    logic [2:0] bit_count_reg, bit_count_next;        // To prevent Latch


    // State Register
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            c_state <= IDLE;
            tx_data_reg <= 8'b0;
            rx_data_reg <= 8'b0;
            sclk_count_reg <= 6'b0;
            bit_count_reg <= 3'b0;
        end else begin
            c_state <= n_state;
            tx_data_reg <= tx_data_next;
            rx_data_reg <= rx_data_next;
            sclk_count_reg <= sclk_count_next;
            bit_count_reg <= bit_count_next;
        end
    end


    // Next State Logic(Combinational) + Output Logic(Combinational)
    always_comb begin
        n_state = c_state;  // �⺻�� ����
        tx_data_next = tx_data_reg;  // �⺻�� ����
        rx_data_next = rx_data_reg;  // �⺻�� ����
        sclk_count_next = sclk_count_reg;  // �⺻�� ����
        bit_count_next = bit_count_reg;  // �⺻�� ����
        tx_ready = 1'b0;  // �⺻�� ����
        done = 1'b0;  // �⺻�� ����
        SCLK = 1'b0;  // CPOL = 0����, �⺻�� ����
        case (c_state)
            IDLE: begin
                    done = 1'b0;          // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                    tx_ready = 1'b1;      // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                    sclk_count_next = 0;
                    bit_count_next = 0;
                if (start) begin
                    n_state = CP0;
                    tx_data_next = tx_data;  //TX data latching
                end else begin
                    n_state = IDLE;
                end
            end
            CP0: begin
                SCLK = 0; // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                if (sclk_count_reg == 49) begin    // Rising Edge
                    rx_data_next = {rx_data[6:0], MISO};  // MSB first ����
                    sclk_count_next = 0;
                    n_state = CP1;
                end else begin
                    sclk_count_next = sclk_count_reg + 1;
                    n_state = CP0;
                end
            end
            CP1: begin
                SCLK = 1; // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                if (sclk_count_reg == 49) begin
                    sclk_count_next = 0;
                    if (bit_count_reg == 7) begin   // Falling Edge
                        bit_count_next = 0;
                        done = 1;
                        n_state = IDLE;
                    end else begin
                        bit_count_next = bit_count_reg + 1;
                        tx_data_next = {tx_data_reg[6:0], 1'b0};  // MSB first ����
                        n_state = CP0;
                    end
                end else begin
                    sclk_count_next = sclk_count_reg + 1;
                    n_state = CP1;
                end
            end
        endcase
    end

    // ��, tx_data, bit_count, sclk_count���� ��ȣ���� ��������ȭ �ߴ°�?
    // => Latch ���� ����.
    // => Combinational logic���� ��ȣ�� ���� ���¸� ������ ��,
    //    �ش� ��ȣ���� ��������ȭ �Ǿ� ���� ������, ��ȣ�� ���� ���¸� �����ϱ� ���� Latch�� ������ �� ����.
    //    �̴� ����ġ ���� ������ �ʷ��� �� ����.
    // ������ ���� �ش� ��ȣ�� Module�� output ��Ʈ���, ��������ȭ ���� �ʾƵ� ��.
    // => Module�� output ��Ʈ�� �⺻������ Combinational logic���� ���� �Ҵ�ޱ� ������,
    //    Latch�� ������ ������ ����. 
    //
    // ��, ����� internal signal���� combinational logic�ӿ��� �� ���� �ٲ�� �ȴٸ�
    // �ش� signal���� ��������ȭ �ؾ���. (LATCH ���� ����)
    // �ݸ鿡, ����� output ��Ʈ���� ��������ȭ ���� �ʾƵ� ��.

    assign MOSI = tx_data_reg[7];  // MSB first ����
    assign rx_data = rx_data_reg;  // ���� ���� ������
endmodule
